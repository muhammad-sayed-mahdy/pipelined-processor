LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

--Instruction Memory
ENTITY rom IS
	GENERIC ( n : integer := 16);
	PORT(
		address : IN  std_logic_vector(10 DOWNTO 0);
		dataout : OUT std_logic_vector(n-1 DOWNTO 0));
END ENTITY rom;

ARCHITECTURE rom_arch OF rom IS

	TYPE rom_type IS ARRAY(0 TO 59) OF std_logic_vector(n-1 DOWNTO 0);
	SIGNAL rom : rom_type := (
		"0000000000000000",
		"0000000000000001",
		"0000000000000010",
		"1100000000000011",
		"1100000000000100",
		"0000000000000101",
		"0000000000000110",
		"0000000000000111",
		"0000000000001000",
		"0000000000001001",
		"0000000000001010",
		"0000000000001011",
		"1100000000001100",
		"0000000000001101",
		"1100100000001110",
		"1100000000001111",
		"0000000000010000",
		"0000000000010001",
		"0000000000010010",
		"0000000000010011",
		"0000000000010100",
		"0000000000010101",
		"0000000000010110",
		"0000000000010111",
		"0000000000011000",
		"0000000000011001",
		"0000000000011010",
		"0000000000011011",
		"0000000000011100",
		"0000000000011101",
		"0000000000011110",
		"0000000000011111",
		"0000000000100000",
		"1100000000100001",
		"1100000000100010",
		"0000000000100011",
		"0000000000100100",
		"0000000000100101",
		"0000000000100110",
		"0000000000100111",
		"0000000000101000",
		"0000000000101001",
		"0000000000101010",
		"0000000000101011",
		"0000000000101100",
		"0000000000101101",
		"0000000000101110",
		"0000000000101111",
		"0000000000110000",
		"0000000000110001",
		"0000000000110010",
		"0000000000110011",
		"0000000000110100",
		"0000000000110101",
		"0000000000110110",
		"0000000000110111",
		"0000000000111000",
		"0000000000111001",
		"0000000000111010",
		"0000000000111011"
	);
	BEGIN
		dataout <= rom(to_integer(unsigned(address)));
END rom_arch;
